library IEEE;
use IEEE.std_logic_1164.all;

package custom_types is
    
    type 2D_matrix is array ( natural range <> ) of std_logic_vector;


end package MIPS_types;